library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity u_rx is
    port (
        clk : in std_logic;
        rst : in std_logic;
        baud_tick_8x : in std_logic;
        rx_i : in std_logic;
        parity_enable : in std_logic;
        parity_even : in std_logic;
        data_bus : out std_logic_vector(7 downto 0);
        LEDR0 : out std_logic;
        data_ready : out std_logic
    );
end entity;

architecture rtl of u_rx is
    component rx_shiftreg is
        port (
            clk : in std_logic;
            rst : in std_logic;
            shift_en : in std_logic;
            rx_bit : in std_logic;
            clear : in std_logic;
            data : out std_logic_vector(7 downto 0)
            --bit_cnt         : out integer range 0 to 7;
            --byte_done       : out std_logic
        );
    end component;

    signal sh_data : std_logic_vector(7 downto 0);

    --Oversampeling signals
    signal bit_cnt : integer range 0 to 7 := 0;
    signal bit_mid_i : std_logic := '0';
    signal shift_en : std_logic;

    -- Signals
    type state_type is (idle, start, data, parity, stop);
    signal state : state_type := idle;
    signal tick_cnt : unsigned(2 downto 0) := (others => '0');
    signal rx_sync : std_logic := '1';
    signal data_ready_i : std_logic := '0';
    signal sh_clear : std_logic := '0';
    signal parity_bit_rx : std_logic := '0';

    -- Main prosess
begin
    -- instans av shiftregisteret
    u_shift : rx_shiftreg
    port map(
        clk => clk,
        rst => rst,
        shift_en => shift_en,
        rx_bit => rx_sync,
        clear => sh_clear,
        data => sh_data
        --bit_cnt         => sh_bit_cnt,
        --byte_done       => sh_byte_done
    );

    process (clk, rst)
    begin
        --Reset logic
        if rst = '1' then
            state <= idle;
            tick_cnt <= (others => '0');
            data_ready_i <= '0';
            rx_sync <= '1';
            shift_en <= '0';
            sh_clear <= '0';

        elsif rising_edge(clk) then
            rx_sync <= rx_i;
            shift_en <= '0';
            data_ready_i <= '0';

            if baud_tick_8x = '1' then
                -- 8x Oversampeling logic
                if tick_cnt = 7 then
                    tick_cnt <= (others => '0');
                else
                    tick_cnt <= tick_cnt + 1;
                end if;

                -- Find middle of bit
                if tick_cnt = 3 then
                    --SHIFTREG_SIGNAL_HERE <= rx_i; -- Stores bit balue
                    bit_mid_i <= '1';
                else
                    bit_mid_i <= '0';
                end if;

                -- UART statemachine logic
                case state is
                    when idle =>
                        sh_clear <= '0';
                        data_ready_i <= '0';
                        tick_cnt <= (others => '0');

                        -- data detected
                        if rx_sync = '0' then
                            state <= start;
                            --initialize counter
                            tick_cnt <= (others => '0');
                        end if;

                    when start =>
                        --sample middle value
                        if tick_cnt = 3 then
                            -- rx line still pulled low
                            if rx_sync = '0' then
                                state <= data;
                            else
                                state <= idle; -- glitch (reset)
                            end if;
                        end if;
                        tick_cnt <= tick_cnt + 1;

                    when data =>
                        if tick_cnt = 3 then
                            shift_en <= '1';

                            if bit_cnt = 7 then
                                bit_cnt <= 0;

                                if parity_enable = '1' then
                                    state <= parity;
                                else
                                    state <= stop;
                                end if;

                            else
                                bit_cnt <= bit_cnt + 1;
                            end if;
                        end if;
                        tick_cnt <= tick_cnt + 1;

                    when parity =>
                        if tick_cnt = 3 then
                            parity_bit_rx <= rx_sync; -- sample received parity bit
                            state <= stop;
                        end if;
                        tick_cnt <= tick_cnt + 1;

                    when stop =>
                        if tick_cnt = 3 then

                            -- STOP bit check
                            if rx_sync = '1' then
                                
                                -- XOR of entire data byte
                                variable p : std_logic := '0';
                            begin
                                for i in 0 to 7 loop
                                    p := p xor sh_data(i);
                                end loop;

                                -- even parity means p must equal received bit
                                -- odd parity means p must NOT equal received bit
                                if parity_enable = '1' then
                                    if parity_even = '1' then
                                        -- EVEN parity
                                        if p = parity_bit_rx then
                                            data_ready_i <= '1';
                                        else
                                            LEDR0 <= '1'; -- parity error
                                        end if;
                                    else
                                        -- ODD parity
                                        if p /= parity_bit_rx then
                                            data_ready_i <= '1';
                                        else
                                            LEDR0 <= '1'; -- parity error
                                        end if;
                                    end if;
                                else
                                    -- parity disabled → always accept data
                                    data_ready_i <= '1';
                                end if;

                                sh_clear <= '1';
                            end if;

                            state <= idle;

                        else
                            tick_cnt <= tick_cnt + 1;
                        end if;
                end case;
            end if;
        end if;
    end process;

    -- separate data-ready process
    process (clk)
    begin
        if rising_edge(clk) then
            if data_ready_i = '1' then
                data_bus <= sh_data;
            elsif baud_tick_8x = '1' then
                data_bus <= (others => '0');
            end if;
        end if;
    end process;

    -- for testbench ?
    bit_mid <= bit_mid_i;

    -- not sure if this is needed
    LEDR0 <= data_ready_i; -- docs just said rx needed a signal to indicate data received
    -- as this one:
    data_ready <= data_ready_i;

    -- this one is implemented as a process now i think
    -- probably ok to delete
    --data_bus    <= (others => '0') when data_ready_i = '0' else sh_data;
end architecture;