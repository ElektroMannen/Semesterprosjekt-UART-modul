library ieee; 
use ieee.std_logic_1164.all;

entity u_baudgen is
	port (
		clk		:	in  std_logic;
		rst_n		:	in  std_logic;
		tick		:	out std_logic
	);
end entity;


architecture rtl of u_baudgen is
begin



end architecture;
