library ieee;
use ieee.std_logic_1164.all;


entity u_ctrl is
	port (
		clk		: in  std_logic;
		rst		: in  std_logic
	);
end entity;


architecture rtl of u_ctrl is

begin
end architecture;
